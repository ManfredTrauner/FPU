`default_nettype none


module tt_um_test1 (
    input  wire [7:0] ui_in,    // Dedicated inputs - connected to the input switches
    output wire [7:0] uo_out,   // Dedicated outputs - connected to the 7 segment display
    input  wire [7:0] uio_in,   // IOs: Bidirectional Input path
    output wire [7:0] uio_out,  // IOs: Bidirectional Output path
    output wire [7:0] uio_oe,   // IOs: Bidirectional Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // will go high when the design is enabled
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);


    // use bidirectionals as outputs
    assign uio_oe = 8'b11111111;
    assign uio_out = 8'hFF;
    assign uo_out = 8'hFF;

    wire reset;
    assign reset = !rst_n;
    
    wire x;
    wire A, B, out1;
    assign x = ui_in[0];
    assign A = ui_in[7];
    assign B = ui_in[6];
    assign out1 = ((~x&A)&A)|(B&x);

    always @(posedge clk or posedge reset) begin
        // if reset, set 
        if (reset) begin
	
        end 
    end
    
    always @(*) begin
//      iresult_mant = operand_a_mant * operand_b_mant;
    end
      


endmodule
